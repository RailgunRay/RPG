    ����          Assembly-CSharp   TestSave+Parametrs   HPxyz       $   }Q&�-��A    