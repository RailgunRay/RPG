    ����          Assembly-CSharp   TestSave+Parametrs   HPxyz       $   ����A    